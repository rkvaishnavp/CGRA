module registers (
    input rs1addr,
    input rs2addr,
    output rs1data,
    output rs2data,
    
    """
    
    """

);
    
endmodule