module cgra_2x2_tb;

